library verilog;
use verilog.vl_types.all;
entity mips32 is
    port(
        CLK             : in     vl_logic
    );
end mips32;
