library verilog;
use verilog.vl_types.all;
entity mips32_testbench is
end mips32_testbench;
